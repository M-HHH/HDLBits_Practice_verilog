module top_module (
    input [7:0] a,
    input [7:0] b,
    output [7:0] s,
    output overflow
); //
 
     assign s = a + b;
    assign overflow = (a[7] == b[7] && a[7] != s[7])?1:0;
    
    //溢出判断方法一 　　用Xf和Yf表示被加数和加数补码的符号位，Zf为补码和的符号位。当出现Xf = Yf= 0两数同为正，而Zf为负,即Zf=1时，有上溢。当出现Xf =Yf = 1两数同为负，而Zf为正，即Zf= 0时，有下溢。 
    //溢出判断方法二 　　当数值最高位有进位位C1=1，符号位没有进位C0=0时，或当数值最高位没有进位位C1=0，符号位有进位C0=1时，结果有溢出。 
    //溢出判断方法三： 用变形补码进行双符号位运算。在变形补码中，正数符号以"00"表示，负数的符号以"11"表示。一般称左边的符号位为第一符号位，右边的符号位为第二符号位。若运算结果的符号位为"01"，则表明有正溢出产生。若运算结果的符号"10"，则表明有负溢出产生。



endmodule
